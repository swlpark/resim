library verilog;
use verilog.vl_types.all;
entity my_region_sv_unit is
end my_region_sv_unit;
