library verilog;
use verilog.vl_types.all;
entity my_solyr_sv_unit is
end my_solyr_sv_unit;
