library verilog;
use verilog.vl_types.all;
entity xbuscore is
    port(
        clk             : in     vl_logic;
        rstn            : in     vl_logic;
        ma0_req         : in     vl_logic;
        xbm0_gnt        : out    vl_logic;
        ma0_select      : in     vl_logic;
        ma0_addr        : in     vl_logic_vector(31 downto 0);
        ma0_data        : in     vl_logic_vector(31 downto 0);
        ma0_rnw         : in     vl_logic;
        ma0_be          : in     vl_logic_vector(3 downto 0);
        xbm0_ack        : out    vl_logic;
        xbm0_data       : out    vl_logic_vector(31 downto 0);
        ma1_req         : in     vl_logic;
        xbm1_gnt        : out    vl_logic;
        ma1_select      : in     vl_logic;
        ma1_addr        : in     vl_logic_vector(31 downto 0);
        ma1_data        : in     vl_logic_vector(31 downto 0);
        ma1_rnw         : in     vl_logic;
        ma1_be          : in     vl_logic_vector(3 downto 0);
        xbm1_ack        : out    vl_logic;
        xbm1_data       : out    vl_logic_vector(31 downto 0);
        ma2_req         : in     vl_logic;
        xbm2_gnt        : out    vl_logic;
        ma2_select      : in     vl_logic;
        ma2_addr        : in     vl_logic_vector(31 downto 0);
        ma2_data        : in     vl_logic_vector(31 downto 0);
        ma2_rnw         : in     vl_logic;
        ma2_be          : in     vl_logic_vector(3 downto 0);
        xbm2_ack        : out    vl_logic;
        xbm2_data       : out    vl_logic_vector(31 downto 0);
        ma3_req         : in     vl_logic;
        xbm3_gnt        : out    vl_logic;
        ma3_select      : in     vl_logic;
        ma3_addr        : in     vl_logic_vector(31 downto 0);
        ma3_data        : in     vl_logic_vector(31 downto 0);
        ma3_rnw         : in     vl_logic;
        ma3_be          : in     vl_logic_vector(3 downto 0);
        xbm3_ack        : out    vl_logic;
        xbm3_data       : out    vl_logic_vector(31 downto 0);
        xbs_select      : out    vl_logic;
        xbs_addr        : out    vl_logic_vector(31 downto 0);
        xbs_data        : out    vl_logic_vector(31 downto 0);
        xbs_rnw         : out    vl_logic;
        xbs_be          : out    vl_logic_vector(3 downto 0);
        sl_ack          : in     vl_logic;
        sl_data         : in     vl_logic_vector(31 downto 0)
    );
end xbuscore;
