library verilog;
use verilog.vl_types.all;
entity error_if is
end error_if;
