library verilog;
use verilog.vl_types.all;
entity my_if is
end my_if;
