library verilog;
use verilog.vl_types.all;
entity null_if is
end null_if;
