library verilog;
use verilog.vl_types.all;
entity icap_virtex_wrapper_sv_unit is
end icap_virtex_wrapper_sv_unit;
